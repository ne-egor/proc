`ifndef __FUNCT_VH
`define __FUNCT_VH

// Здесь хранятся макроопределения для кодов арифметико-логических операций модельной архитектуры.
// Названия говорят сами за себя.
`define FUNCT_ADD  4'b1000
`define FUNCT_SUB  4'b1010
`define FUNCT_AND  4'b0100
`define FUNCT_OR   4'b0110
`define FUNCT_SLTU 4'b0010
`define FUNCT_SLT  4'b0011

`endif // __FUNCT_VH
